

library IEEE;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.STD_LOGIC_1164.all;



entity MemDOs is port(
	clk: 			in std_logic; 			 
	Write_Dat : 	in STD_LOGIC_VECTOR(63 downto 0);
	W_Enable: 		in std_logic; 	
	Adress: 		in std_logic_vector(7 downto 0);	
--	Read: 			in std_logic;
	Read_Dat: 		out std_logic_vector(63 downto 0)
	);
end MemDOs;



architecture MemDOs of MemDOs is
type Dato_Mem2 is array (0 to 255) of std_logic_vector(63 downto 0);
signal Dato : Dato_Mem2 :=(	 

	x"0000000000000001",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"0000000000000023",x"0000000000000041",
	x"0000000000000015",x"0000000000000000",x"0000000000000030",x"000000000000000f",

	x"0000000000000010",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f",	
	
	x"0000000000000020",x"0000000000000021",x"0000000000000034",x"0000000000000023",
	x"0000000000000024",x"0000000000000025",x"0000000000000026",x"0000000000000027",
	x"0000000000000028",x"0000000000000029",x"000000000000002a",x"000000000000002b",
	x"000000000000002c",x"000000000000002d",x"000000000000002e",x"000000000000002f",

	x"0000000000000030",x"0000000000000000",x"0000000000000032",x"0000000000000033",
	x"0000000000000034",x"0000000000000035",x"0000000000000036",x"0000000000000037",
	x"0000000000000038",x"0000000000000039",x"000000000000003a",x"000000000000003b",
	x"000000000000003c",x"000000000000003d",x"000000000000003e",x"000000000000003f",
	
	x"0000000000000000",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"0000000000000000",

	x"0000000000000050",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000039",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000000f",	
	
	x"000000000000005f",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000000",
	x"000000000000006f",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"0000000000000000",

	x"000000000000007f",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f",  
	
	x"0000000000000000",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"000000000000000f",

	x"0000000000000010",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f",	
	
	x"0000000000000000",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"000000000000000f",

	x"0000000000000010",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f",
	
	x"0000000000000000",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"000000000000000f",

	x"0000000000000010",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f",	
	
	x"0000000000000000",x"0000000000000001",x"0000000000000002",x"0000000000000003",
	x"0000000000000004",x"0000000000000005",x"0000000000000006",x"0000000000000007",
	x"0000000000000008",x"0000000000000009",x"000000000000000a",x"000000000000000b",
	x"000000000000000c",x"000000000000000d",x"000000000000000e",x"000000000000000f",

	x"0000000000000010",x"0000000000000011",x"0000000000000012",x"0000000000000013",
	x"0000000000000014",x"0000000000000015",x"0000000000000016",x"0000000000000017",
	x"0000000000000018",x"0000000000000019",x"000000000000001a",x"000000000000001b",
	x"000000000000001c",x"000000000000001d",x"000000000000001e",x"000000000000001f"

);
begin
	process	(clk,Adress,Write_Dat,W_Enable)
		begin
			if (W_Enable = '1' and rising_edge(clk)) then
				Dato(conv_integer(Adress(7 downto 0)))	<= Write_Dat;
			end if;
			
			Read_Dat	<= Dato(conv_integer(Adress (7 downto 0)));	
	end process;

end MemDOs;
